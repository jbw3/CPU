// Decoder5to32
// John Wilkes

module Decoder5to32(input [4:0] I, output reg [31:0] O);

    always @(I)
        case(I)
             0: O <= 32'h00000001;
             1: O <= 32'h00000002;
             2: O <= 32'h00000004;
             3: O <= 32'h00000008;
             4: O <= 32'h00000010;
             5: O <= 32'h00000020;
             6: O <= 32'h00000040;
             7: O <= 32'h00000080;
             8: O <= 32'h00000100;
             9: O <= 32'h00000200;
            10: O <= 32'h00000400;
            11: O <= 32'h00000800;
            12: O <= 32'h00001000;
            13: O <= 32'h00002000;
            14: O <= 32'h00004000;
            15: O <= 32'h00008000;
            16: O <= 32'h00010000;
            17: O <= 32'h00020000;
            18: O <= 32'h00040000;
            19: O <= 32'h00080000;
            20: O <= 32'h00100000;
            21: O <= 32'h00200000;
            22: O <= 32'h00400000;
            23: O <= 32'h00800000;
            24: O <= 32'h01000000;
            25: O <= 32'h02000000;
            26: O <= 32'h04000000;
            27: O <= 32'h08000000;
            28: O <= 32'h10000000;
            29: O <= 32'h20000000;
            30: O <= 32'h40000000;
            31: O <= 32'h80000000;
        endcase

endmodule
